* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT fig3_1layout Vdd A B C D Y gnd
** N=10 EP=7 IP=0 FDC=8
M0 Y A gnd gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=1025 $Y=-785 $D=0
M1 4 B Y gnd N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=3655 $Y=-785 $D=0
M2 gnd C 4 gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=4345 $Y=-785 $D=0
M3 gnd D Y gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=6425 $Y=-785 $D=0
M4 5 A Vdd Vdd P_18 L=1.8e-07 W=3e-06 AD=7.65e-13 AS=1.47e-12 PD=5.1e-07 PS=3.98e-06 $X=1025 $Y=5330 $D=1
M5 8 B 5 Vdd P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=7.65e-13 PD=3.98e-06 PS=5.1e-07 $X=1715 $Y=5330 $D=1
M6 8 C 5 Vdd P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06 $X=4345 $Y=5330 $D=1
M7 Y D 8 Vdd P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06 $X=6425 $Y=5330 $D=1
.ENDS
***************************************
