/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2022 Spring ---------------------- //
// ---------------------- Version : v.1.10  ---------------------- //
// ---------------------- Date : 2022.04.13 ---------------------- //
// ------------------------- USS module ---------------------------//
// ----------------- Feb. 2022 Willie authored --------------------//
/////////////////////////////////////////////////////////////////////

module USS(clk, rst, X_in, X_c, Y_c, neighbor_sel);

// ---------------------- input  ---------------------- //
	input clk;
	input rst;
	input [2:0] X_in;
	input [2:0] X_c;
	input [2:0] Y_c;
	
// ---------------------- output  ---------------------- //
	output [15:0] neighbor_sel;
	
// ---------------------- Write down Your design below  ---------------------- //


endmodule

