* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT fig2_2layout Clk D Q Vdd gnd
** N=12 EP=5 IP=0 FDC=20
M0 2 Clk gnd gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=3205 $Y=3510 $D=0
M1 4 2 D gnd N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=6060 $Y=3510 $D=0
M2 5 Clk 4 gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=6750 $Y=3510 $D=0
M3 gnd 6 5 gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=8970 $Y=3510 $D=0
M4 gnd 4 6 gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=12060 $Y=3510 $D=0
M5 7 Clk gnd gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=14725 $Y=3510 $D=0
M6 8 Clk 6 gnd N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17580 $Y=3510 $D=0
M7 9 7 8 gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=18270 $Y=3510 $D=0
M8 gnd Q 9 gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=20490 $Y=3510 $D=0
M9 gnd 8 Q gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=22705 $Y=3510 $D=0
M10 2 Clk Vdd Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06 $X=3205 $Y=8335 $D=1
M11 4 Clk D Vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=6060 $Y=8335 $D=1
M12 5 2 4 Vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=6750 $Y=8335 $D=1
M13 Vdd 6 5 Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06 $X=8970 $Y=8335 $D=1
M14 Vdd 4 6 Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06 $X=12060 $Y=8335 $D=1
M15 7 Clk Vdd Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06 $X=14725 $Y=8335 $D=1
M16 8 7 6 Vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17580 $Y=8335 $D=1
M17 9 Clk 8 Vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=18270 $Y=8335 $D=1
M18 Vdd Q 9 Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06 $X=20490 $Y=8335 $D=1
M19 Vdd 8 Q Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06 $X=22705 $Y=8335 $D=1
.ENDS
***************************************
