* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT hw3_2b Vin gnd Vdd
** N=7 EP=3 IP=0 FDC=10
M0 2 Vin gnd gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=150 $Y=2455 $D=0
M1 3 2 gnd gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=2085 $Y=2455 $D=0
M2 4 3 gnd gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=3925 $Y=2455 $D=0
M3 5 4 gnd gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=5870 $Y=2455 $D=0
M4 Vin 5 gnd gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=7845 $Y=2455 $D=0
M5 2 Vin Vdd Vdd P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06 $X=150 $Y=7870 $D=1
M6 3 2 Vdd Vdd P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06 $X=2085 $Y=7870 $D=1
M7 4 3 Vdd Vdd P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06 $X=3925 $Y=7870 $D=1
M8 5 4 Vdd Vdd P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06 $X=5870 $Y=7870 $D=1
M9 Vin 5 Vdd Vdd P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06 $X=7845 $Y=7870 $D=1
.ENDS
***************************************
