************************************************************************
* auCdl Netlist:
* 
* Library Name:  Pb1
* Top Cell Name: fig3_1
* View Name:     schematic
* Netlisted on:  Mar 17 20:38:08 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: Pb1
* Cell Name:    fig3_1
* View Name:    schematic
************************************************************************

.SUBCKT fig3_1 A B C D Vdd Y gnd
*.PININFO A:I B:I C:I D:I Vdd:I gnd:I Y:O
MM3 Y D gnd gnd N_18 W=1u L=180n
MM2 net25 C gnd gnd N_18 W=1u L=180n
MM1 Y B net25 gnd N_18 W=1u L=180n
MM0 Y A gnd gnd N_18 W=1u L=180n
MM5 Y D net20 Vdd P_18 W=3u L=180n
MM6 net20 C net21 Vdd P_18 W=3u L=180n
MM4 net20 B net21 Vdd P_18 W=3u L=180n
MM7 net21 A Vdd Vdd P_18 W=3u L=180n
.ENDS

