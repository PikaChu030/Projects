* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT fig3_2layout A B Vdd C gnd Y
** N=8 EP=6 IP=0 FDC=6
M0 2 A gnd gnd N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=610 $Y=-295 $D=0
M1 Y B 2 gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=1300 $Y=-295 $D=0
M2 gnd C Y gnd N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=3380 $Y=-295 $D=0
M3 6 A Vdd Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06 $X=610 $Y=4780 $D=1
M4 6 B Vdd Vdd P_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06 $X=2690 $Y=4780 $D=1
M5 Y C 6 Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=3380 $Y=4780 $D=1
.ENDS
***************************************
