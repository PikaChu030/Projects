* SPICE NETLIST
***************************************

.SUBCKT RM1 A B
.ENDS
***************************************
.SUBCKT RM2 A B
.ENDS
***************************************
.SUBCKT RM3 A B
.ENDS
***************************************
.SUBCKT RM4 A B
.ENDS
***************************************
.SUBCKT RM5 A B
.ENDS
***************************************
.SUBCKT RM6 A B
.ENDS
***************************************
.SUBCKT DN A B
.ENDS
***************************************
.SUBCKT DP A B
.ENDS
***************************************
.SUBCKT L_SLCR20K_RF POS NEG SUB
.ENDS
***************************************
.SUBCKT PAD_RF POS NEG
.ENDS
***************************************
.SUBCKT Nand B GND OUT A VDD
** N=6 EP=5 IP=0 FDC=4
M0 GND B 4 GND N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.525e-13 PD=1.52e-06 PS=1.51e-06 $X=-2470 $Y=-2940 $D=0
M1 4 A OUT GND N_18 L=1.8e-07 W=5e-07 AD=2.5e-13 AS=2.45e-13 PD=1.5e-06 PS=1.48e-06 $X=1385 $Y=-2940 $D=0
M2 OUT B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=5e-13 AS=4.9e-13 PD=2e-06 PS=1.98e-06 $X=-2465 $Y=-440 $D=1
M3 VDD A OUT VDD P_18 L=1.8e-07 W=1e-06 AD=5.3e-13 AS=4.9e-13 PD=2.06e-06 PS=1.98e-06 $X=1385 $Y=-440 $D=1
.ENDS
***************************************
