/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2022 Spring ---------------------- //
// ---------------------- Version : v.1.10  ---------------------- //
// ---------------------- Date : 2022.04.13 ---------------------- //
// ------------------------ VEP module --------------------------//
// ----------------- Feb. 2022 Willie authored --------------------//
/////////////////////////////////////////////////////////////////////

module VEP(clk, rst, W_update, D_update, neighbor_sel, pixel,
				d0, d1, d2, d3, d4, d5, d6, d7, w0, w1, w2, w3, w4, w5, w6, w7);

// ---------------------- input  ---------------------- //
	input clk; 
	input rst; 
	input W_update;
	input D_update;
	input [15:0] neighbor_sel; 
	input [23:0] pixel; 
	
// ---------------------- output  ---------------------- //
	output [10:0] d0;
	output [10:0] d1;
	output [10:0] d2;
	output [10:0] d3;
	output [10:0] d4;
	output [10:0] d5;
	output [10:0] d6;
	output [10:0] d7;
	output [23:0] w0;
	output [23:0] w1;
	output [23:0] w2;
	output [23:0] w3;
	output [23:0] w4;
	output [23:0] w5;
	output [23:0] w6;
	output [23:0] w7;
	
// ---------------------- Write down Your design below  ---------------------- //


endmodule
