************************************************************************
* auCdl Netlist:
* 
* Library Name:  Pb1
* Top Cell Name: INV
* View Name:     schematic
* Netlisted on:  Apr 12 21:43:12 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: Pb1
* Cell Name:    INV
* View Name:    schematic
************************************************************************

.SUBCKT INV Vdd gnd in out
*.PININFO Vdd:I gnd:I in:I out:O
MMN2 out in gnd gnd N_18 W=2u L=180.00n
MMN1 out in Vdd Vdd P_18 W=6u L=180n
.ENDS

