/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2022 Spring ---------------------- //
// ---------------------- Editor : JulianaLu --------------------- //
// ---------------------- Version : v.1.00  ---------------------- //
// ---------------------- Date : 2022.02.15 ---------------------- //
// ----------------------    Manhattan      ---------------------- //
/////////////////////////////////////////////////////////////////////

`timescale 1ns/10ps
`define RGB_DataSize 24
`define D_DataSize 10
// ---------------------- define ---------------------- //

module Manhattan(clk,
                 rst,
                 clear,
                 c_en,
                 if_en,
                 c_in0,
                 c_in1,
                 c_in2,
                 c_in3,
                 c_in4,
                 c_in5,
                 c_in6,
                 c_in7,
                 if_in,
                 d_0,
                 d_1,
                 d_2,
                 d_3,
                 d_4,
                 d_5,
                 d_6,
                 d_7);

  // ---------------------- input  ---------------------- //
  input  clk;
  input  rst;
  input  clear;
  input  c_en;
  input  if_en;
  input   [`RGB_DataSize-1:0] c_in0, c_in1, c_in2, c_in3, c_in4, c_in5, c_in6, c_in7;
  input   [`RGB_DataSize-1:0] if_in;

  // ---------------------- output ---------------------- //
  output  [`D_DataSize-1:0] d_0, d_1, d_2, d_3, d_4, d_5, d_6, d_7;

  // ---------------------- Write down Your design below  ---------------------- //
  reg  [`RGB_DataSize-1:0] t_0,t_1,t_2,t_3,t_4,t_5,t_6,t_7;
  reg  [`RGB_DataSize-1:0] t_in;

  always @(posedge clk or rst) begin
          if (rst == 1'b1) begin
                  t_0 <=24'b0;
                  t_1 <=24'b0;
                  t_2 <=24'b0;
                  t_3 <=24'b0;
                  t_4 <=24'b0;
                  t_5 <=24'b0;
                  t_6 <=24'b0;
                  t_7 <=24'b0;
                  t_in<=24'b0;
          end
          else begin
                  if (clear == 1'b1) begin
                        t_0 <=24'b0;
                        t_1 <=24'b0;
                        t_2 <=24'b0;
                        t_3 <=24'b0;
                        t_4 <=24'b0;
                        t_5 <=24'b0;
                        t_6 <=24'b0;
                        t_7 <=24'b0;
                        t_in<=24'b0;
                  end
                  else begin
                          if(c_en == 1'b1)begin
                                  t_0 <= c_in0;
                                  t_1 <= c_in1;
                                  t_2 <= c_in2;
                                  t_3 <= c_in3;
                                  t_4 <= c_in4;
                                  t_5 <= c_in5;
                                  t_6 <= c_in6;
                                  t_7 <= c_in7;
                          end
                          if(if_en == 1'b1)begin
                                  t_in <= if_in;
                          end 
                  end
          end
  end
      assign d_0 = ((t_in[7:0] >= t_0[7:0])?t_in[7:0] - t_0[7:0] : t_0[7:0] - t_in[7:0] ) + 
                   ((t_in[15:8] >= t_0[15:8])?t_in[15:8] - t_0[15:8] : t_0[15:8] - t_in[15:8] ) +
                   ((t_in[23:16] >= t_0[23:16])?t_in[23:16] - t_0[23:16] : t_0[23:16] - t_in[23:16] );

      assign d_1 = ((t_in[7:0] >= t_1[7:0])?t_in[7:0] - t_1[7:0] : t_1[7:0] - t_in[7:0] ) + 
                   ((t_in[15:8] >= t_1[15:8])?t_in[15:8] - t_1[15:8] : t_1[15:8] - t_in[15:8] ) +
                   ((t_in[23:16] >= t_1[23:16])?t_in[23:16] - t_1[23:16] : t_1[23:16] - t_in[23:16] );

      assign d_2 = ((t_in[7:0] >= t_1[7:0])?t_in[7:0] - t_2[7:0] : t_2[7:0] - t_in[7:0] ) + 
                   ((t_in[15:8] >= t_2[15:8])?t_in[15:8] - t_2[15:8] : t_2[15:8] - t_in[15:8] ) +
                   ((t_in[23:16] >= t_2[23:16])?t_in[23:16] - t_2[23:16] : t_2[23:16] - t_in[23:16] );

      assign d_3 = ((t_in[7:0] >= t_3[7:0])?t_in[7:0] - t_3[7:0] : t_3[7:0] - t_in[7:0] ) + 
                   ((t_in[15:8] >= t_3[15:8])?t_in[15:8] - t_3[15:8] : t_3[15:8] - t_in[15:8] ) +
                   ((t_in[23:16] >= t_3[23:16])?t_in[23:16] - t_3[23:16] : t_3[23:16] - t_in[23:16] );

      assign d_4 = ((t_in[7:0] >= t_4[7:0])?t_in[7:0] - t_4[7:0] : t_4[7:0] - t_in[7:0] ) + 
                   ((t_in[15:8] >= t_4[15:8])?t_in[15:8] - t_4[15:8] : t_4[15:8] - t_in[15:8] ) +
                   ((t_in[23:16] >= t_4[23:16])?t_in[23:16] - t_4[23:16] : t_4[23:16] - t_in[23:16] );

      assign d_5 = ((t_in[7:0] >= t_5[7:0])?t_in[7:0] - t_5[7:0] : t_5[7:0] - t_in[7:0] ) + 
                   ((t_in[15:8] >= t_5[15:8])?t_in[15:8] - t_5[15:8] : t_5[15:8] - t_in[15:8] ) +
                   ((t_in[23:16] >= t_5[23:16])?t_in[23:16] - t_5[23:16] : t_5[23:16] - t_in[23:16] );

      assign d_6 = ((t_in[7:0] >= t_6[7:0])?t_in[7:0] - t_6[7:0] : t_6[7:0] - t_in[7:0] ) + 
                   ((t_in[15:8] >= t_6[15:8])?t_in[15:8] - t_6[15:8] : t_6[15:8] - t_in[15:8] ) +
                   ((t_in[23:16] >= t_6[23:16])?t_in[23:16] - t_6[23:16] : t_6[23:16] - t_in[23:16] );

      assign d_7 = ((t_in[7:0] >= t_7[7:0])?t_in[7:0] - t_7[7:0] : t_7[7:0] - t_in[7:0] ) + 
                   ((t_in[15:8] >= t_7[15:8])?t_in[15:8] - t_7[15:8] : t_7[15:8] - t_in[15:8] ) +
                   ((t_in[23:16] >= t_7[23:16])?t_in[23:16] - t_7[23:16] : t_7[23:16] - t_in[23:16] );
  endmodule
