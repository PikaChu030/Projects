* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT fig1_6layout D0 Y D1 S gnd Vdd
** N=7 EP=6 IP=0 FDC=6
M0 Y 4 D0 gnd N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=2.89e-12 PD=5.1e-07 PS=4.89e-06 $X=8155 $Y=-5340 $D=0
M1 D1 S Y gnd N_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=8845 $Y=-5340 $D=0
M2 gnd S 4 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=4.9e-13 PD=1.48e-06 PS=2.46e-06 $X=11585 $Y=-5340 $D=0
M3 Y S D0 Vdd P_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=2.89e-12 PD=5.1e-07 PS=4.89e-06 $X=8155 $Y=1625 $D=1
M4 D1 4 Y Vdd P_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=8845 $Y=1625 $D=1
M5 Vdd S 4 Vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=9.8e-13 PD=1.98e-06 PS=2.96e-06 $X=11585 $Y=1735 $D=1
.ENDS
***************************************
